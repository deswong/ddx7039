#
#   flash_edb9312_ken.cdl
# 
#   FLASH memory - Hardware support on kenwood board
#   data 2006.06.05

#====================================================================
#
#      flash_edb9312.cdl
#
#      FLASH memory - Hardware support on Cirrus Logic EP93xx eval board
#
#====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
#-------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.
# All Rights Reserved.                                                     
#-------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas, hmt
# Original data:  gthomas
# Contributors:   gthomas
# Date:           2001-04-23
#
#####DESCRIPTIONEND####
#
#====================================================================

cdl_package CYGPKG_DEVS_FLASH_EDB9312_KEN {
    display       "Cirrus Logic EP93xx (EDB9312) FLASH memory support"
    description   "FLASH memory device support for Cirrus Logic EDB9312"

    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH
    requires	  CYGPKG_HAL_ARM_ARM9_EP93XX

    implements    CYGHWR_IO_FLASH_DEVICE

    compile       edb9312_flash.c


    # Arguably this should do in the generic package
    # but then there is a logic loop so you can never enable it.
    cdl_interface CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED {
        display   "Generic AMD FLASH driver required"
    }

    implements    CYGINT_DEVS_FLASH_AMD_AM29XXXXX_REQUIRED
    requires      CYGHWR_DEVS_FLASH_AMD_S29GL256N
    requires      CYGHWR_DEVS_FLASH_AMD_S29GL128N
    requires      CYGHWR_DEVS_FLASH_AMD_S29PL127J
}
